-- Test File --